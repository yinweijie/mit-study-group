import ProcTypes::*;
import MemTypes::*;
import Types::*;
import CacheTypes::*;
import MessageFifo::*;
import Vector::*;

module mkPPP(MessageGet c2m, MessagePut m2c, WideMem mem, Empty ifc);
    // TODO: Exercise 4
endmodule
