import Ehr::*;
import Vector::*;
import FIFO::*;

interface Fifo#(numeric type n, type t);
    method Action enq(t x);
    method Action deq;
    method t first;
    method Bool notEmpty;
endinterface

module mkFifo(Fifo#(3, t)) provisos (Bits#(t, tSz));
    // TODO: Exercise 1
    method Action enq(t x);
    endmethod

    method Action deq;
    endmethod

    method t first;
        return ?;
    endmethod

    method Bool notEmpty;
        return False;
    endmethod
endmodule

// Two elements conflict-free FIFO given as black box
module mkCFFifo(Fifo#(2, t)) provisos (Bits#(t, tSz));
    Ehr#(2, t) da <- mkEhr(?);
    Ehr#(2, Bool) va <- mkEhr(False);
    Ehr#(2, t) db <- mkEhr(?);
    Ehr#(2, Bool) vb <- mkEhr(False);

    rule canonicalize;
        if (vb[1] && !va[1]) begin
            da[1] <= db[1];
            va[1] <= True;
            vb[1] <= False;
        end
    endrule

    method Action enq(t x) if (!vb[0]);
        db[0] <= x;
        vb[0] <= True;
    endmethod

    method Action deq if (va[0]);
        va[0] <= False;
    endmethod

    method t first if (va[0]);
        return da[0];
    endmethod

    method Bool notEmpty;
        return va[0];
    endmethod
endmodule

module mkCF3Fifo(Fifo#(3, t)) provisos (Bits#(t, tSz));
    // TODO: optional helper FIFO
    method Action enq(t x);
    endmethod

    method Action deq;
    endmethod

    method t first;
        return ?;
    endmethod

    method Bool notEmpty;
        return False;
    endmethod
endmodule
